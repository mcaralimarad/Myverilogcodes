    module not_my(a,b);//Not gate
    input a;
    output b;
    assign b = ~a;
    endmodule
