module muxprimitive (F, A, I0, I1);
output F;
input A, I0, I1; 

mux1(F, A, I0, I1);

endmodule