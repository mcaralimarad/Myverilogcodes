module and_my(a,b,c); //and gate
    input a,b;
    output c;
    assign c =  a & b;
    endmodule
