    module or_my(a,b,c); //or gate
    input a,b;
    output c;
    assign c =  a || b;
    endmodule
